
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.echo_pkg.ALL;

ENTITY flanger IS
  PORT( clk                               :   IN    std_logic;
        reset                             :   IN    std_logic;
        clk_enable                        :   IN    std_logic;
        In1                               :   IN    std_logic_vector(7 DOWNTO 0);  -- int8
        ce_out                            :   OUT   std_logic;
        Out1                              :   OUT   std_logic_vector(7 DOWNTO 0)  -- int8
        );
END flanger;


ARCHITECTURE rtl OF flanger IS

  -- Signals
  SIGNAL enb                              : std_logic;
  SIGNAL In1_signed                       : signed(7 DOWNTO 0);  -- int8
  SIGNAL Delay_reg                        : vector_of_signed8(0 TO 479);  -- sfix8 [6000]
  SIGNAL Delay_out1                       : signed(7 DOWNTO 0);  -- int8
  SIGNAL attenuation_cast                 : signed(15 DOWNTO 0);  -- sfix16_En7
  SIGNAL attenuation_out1                 : signed(7 DOWNTO 0);  -- int8
  SIGNAL attenuation_cast2                 : signed(15 DOWNTO 0);  -- sfix16_En7
  SIGNAL attenuation_out2                 : signed(7 DOWNTO 0);  -- int8
  SIGNAL Sum_out1                         : signed(7 DOWNTO 0);  -- int8
  SIGNAL sin_pos											: INTEGER RANGE 0 TO 480;

BEGIN
  In1_signed <= signed(In1);

  enb <= clk_enable;

  Delay_process : PROCESS (clk, reset)
  VARIABLE count1  :  INTEGER RANGE 0 TO 150 := 0;  --timing for clock generation
  VARIABLE count2  :  INTEGER RANGE 0 TO 480 := 0;
  BEGIN
    IF reset = '1' THEN
      Delay_reg <= (OTHERS => to_signed(16#00#, 8));
    ELSIF clk'EVENT AND clk = '1' THEN
      IF enb = '1' THEN
			IF(count1 < 150) THEN
				count1 := count1 + 1;
			ELSE
				count1 := 0;
				IF(count2 < 480) THEN
					count2 := count2 + 1;
				ELSE
					count2 := 0;
				END IF;
			END IF;
			CASE count2 IS
				WHEN  0  =>
					 sin_pos <= 0 ;
				WHEN  1  =>
					 sin_pos <= 0 ;
				WHEN  2  =>
					 sin_pos <= 0 ;
				WHEN  3  =>
					 sin_pos <= 0 ;
				WHEN  4  =>
					 sin_pos <= 0 ;
				WHEN  5  =>
					 sin_pos <= 0 ;
				WHEN  6  =>
					 sin_pos <= 0 ;
				WHEN  7  =>
					 sin_pos <= 1 ;
				WHEN  8  =>
					 sin_pos <= 1 ;
				WHEN  9  =>
					 sin_pos <= 1 ;
				WHEN  10  =>
					 sin_pos <= 2 ;
				WHEN  11  =>
					 sin_pos <= 2 ;
				WHEN  12  =>
					 sin_pos <= 2 ;
				WHEN  13  =>
					 sin_pos <= 3 ;
				WHEN  14  =>
					 sin_pos <= 4 ;
				WHEN  15  =>
					 sin_pos <= 4 ;
				WHEN  16  =>
					 sin_pos <= 5 ;
				WHEN  17  =>
					 sin_pos <= 5 ;
				WHEN  18  =>
					 sin_pos <= 6 ;
				WHEN  19  =>
					 sin_pos <= 7 ;
				WHEN  20  =>
					 sin_pos <= 8 ;
				WHEN  21  =>
					 sin_pos <= 9 ;
				WHEN  22  =>
					 sin_pos <= 9 ;
				WHEN  23  =>
					 sin_pos <= 10 ;
				WHEN  24  =>
					 sin_pos <= 11 ;
				WHEN  25  =>
					 sin_pos <= 12 ;
				WHEN  26  =>
					 sin_pos <= 13 ;
				WHEN  27  =>
					 sin_pos <= 14 ;
				WHEN  28  =>
					 sin_pos <= 15 ;
				WHEN  29  =>
					 sin_pos <= 17 ;
				WHEN  30  =>
					 sin_pos <= 18 ;
				WHEN  31  =>
					 sin_pos <= 19 ;
				WHEN  32  =>
					 sin_pos <= 20 ;
				WHEN  33  =>
					 sin_pos <= 22 ;
				WHEN  34  =>
					 sin_pos <= 23 ;
				WHEN  35  =>
					 sin_pos <= 24 ;
				WHEN  36  =>
					 sin_pos <= 26 ;
				WHEN  37  =>
					 sin_pos <= 27 ;
				WHEN  38  =>
					 sin_pos <= 29 ;
				WHEN  39  =>
					 sin_pos <= 30 ;
				WHEN  40  =>
					 sin_pos <= 32 ;
				WHEN  41  =>
					 sin_pos <= 33 ;
				WHEN  42  =>
					 sin_pos <= 35 ;
				WHEN  43  =>
					 sin_pos <= 37 ;
				WHEN  44  =>
					 sin_pos <= 38 ;
				WHEN  45  =>
					 sin_pos <= 40 ;
				WHEN  46  =>
					 sin_pos <= 42 ;
				WHEN  47  =>
					 sin_pos <= 44 ;
				WHEN  48  =>
					 sin_pos <= 45 ;
				WHEN  49  =>
					 sin_pos <= 47 ;
				WHEN  50  =>
					 sin_pos <= 49 ;
				WHEN  51  =>
					 sin_pos <= 51 ;
				WHEN  52  =>
					 sin_pos <= 53 ;
				WHEN  53  =>
					 sin_pos <= 55 ;
				WHEN  54  =>
					 sin_pos <= 57 ;
				WHEN  55  =>
					 sin_pos <= 59 ;
				WHEN  56  =>
					 sin_pos <= 61 ;
				WHEN  57  =>
					 sin_pos <= 63 ;
				WHEN  58  =>
					 sin_pos <= 65 ;
				WHEN  59  =>
					 sin_pos <= 68 ;
				WHEN  60  =>
					 sin_pos <= 70 ;
				WHEN  61  =>
					 sin_pos <= 72 ;
				WHEN  62  =>
					 sin_pos <= 74 ;
				WHEN  63  =>
					 sin_pos <= 77 ;
				WHEN  64  =>
					 sin_pos <= 79 ;
				WHEN  65  =>
					 sin_pos <= 81 ;
				WHEN  66  =>
					 sin_pos <= 84 ;
				WHEN  67  =>
					 sin_pos <= 86 ;
				WHEN  68  =>
					 sin_pos <= 88 ;
				WHEN  69  =>
					 sin_pos <= 91 ;
				WHEN  70  =>
					 sin_pos <= 93 ;
				WHEN  71  =>
					 sin_pos <= 96 ;
				WHEN  72  =>
					 sin_pos <= 98 ;
				WHEN  73  =>
					 sin_pos <= 101 ;
				WHEN  74  =>
					 sin_pos <= 104 ;
				WHEN  75  =>
					 sin_pos <= 106 ;
				WHEN  76  =>
					 sin_pos <= 109 ;
				WHEN  77  =>
					 sin_pos <= 111 ;
				WHEN  78  =>
					 sin_pos <= 114 ;
				WHEN  79  =>
					 sin_pos <= 117 ;
				WHEN  80  =>
					 sin_pos <= 119 ;
				WHEN  81  =>
					 sin_pos <= 122 ;
				WHEN  82  =>
					 sin_pos <= 125 ;
				WHEN  83  =>
					 sin_pos <= 128 ;
				WHEN  84  =>
					 sin_pos <= 131 ;
				WHEN  85  =>
					 sin_pos <= 133 ;
				WHEN  86  =>
					 sin_pos <= 136 ;
				WHEN  87  =>
					 sin_pos <= 139 ;
				WHEN  88  =>
					 sin_pos <= 142 ;
				WHEN  89  =>
					 sin_pos <= 145 ;
				WHEN  90  =>
					 sin_pos <= 148 ;
				WHEN  91  =>
					 sin_pos <= 151 ;
				WHEN  92  =>
					 sin_pos <= 153 ;
				WHEN  93  =>
					 sin_pos <= 156 ;
				WHEN  94  =>
					 sin_pos <= 159 ;
				WHEN  95  =>
					 sin_pos <= 162 ;
				WHEN  96  =>
					 sin_pos <= 165 ;
				WHEN  97  =>
					 sin_pos <= 168 ;
				WHEN  98  =>
					 sin_pos <= 171 ;
				WHEN  99  =>
					 sin_pos <= 174 ;
				WHEN  100  =>
					 sin_pos <= 177 ;
				WHEN  101  =>
					 sin_pos <= 180 ;
				WHEN  102  =>
					 sin_pos <= 183 ;
				WHEN  103  =>
					 sin_pos <= 187 ;
				WHEN  104  =>
					 sin_pos <= 190 ;
				WHEN  105  =>
					 sin_pos <= 193 ;
				WHEN  106  =>
					 sin_pos <= 196 ;
				WHEN  107  =>
					 sin_pos <= 199 ;
				WHEN  108  =>
					 sin_pos <= 202 ;
				WHEN  109  =>
					 sin_pos <= 205 ;
				WHEN  110  =>
					 sin_pos <= 208 ;
				WHEN  111  =>
					 sin_pos <= 211 ;
				WHEN  112  =>
					 sin_pos <= 214 ;
				WHEN  113  =>
					 sin_pos <= 218 ;
				WHEN  114  =>
					 sin_pos <= 221 ;
				WHEN  115  =>
					 sin_pos <= 224 ;
				WHEN  116  =>
					 sin_pos <= 227 ;
				WHEN  117  =>
					 sin_pos <= 230 ;
				WHEN  118  =>
					 sin_pos <= 233 ;
				WHEN  119  =>
					 sin_pos <= 236 ;
				WHEN  120  =>
					 sin_pos <= 239 ;
				WHEN  121  =>
					 sin_pos <= 243 ;
				WHEN  122  =>
					 sin_pos <= 246 ;
				WHEN  123  =>
					 sin_pos <= 249 ;
				WHEN  124  =>
					 sin_pos <= 252 ;
				WHEN  125  =>
					 sin_pos <= 255 ;
				WHEN  126  =>
					 sin_pos <= 258 ;
				WHEN  127  =>
					 sin_pos <= 261 ;
				WHEN  128  =>
					 sin_pos <= 265 ;
				WHEN  129  =>
					 sin_pos <= 268 ;
				WHEN  130  =>
					 sin_pos <= 271 ;
				WHEN  131  =>
					 sin_pos <= 274 ;
				WHEN  132  =>
					 sin_pos <= 277 ;
				WHEN  133  =>
					 sin_pos <= 280 ;
				WHEN  134  =>
					 sin_pos <= 283 ;
				WHEN  135  =>
					 sin_pos <= 286 ;
				WHEN  136  =>
					 sin_pos <= 289 ;
				WHEN  137  =>
					 sin_pos <= 292 ;
				WHEN  138  =>
					 sin_pos <= 296 ;
				WHEN  139  =>
					 sin_pos <= 299 ;
				WHEN  140  =>
					 sin_pos <= 302 ;
				WHEN  141  =>
					 sin_pos <= 305 ;
				WHEN  142  =>
					 sin_pos <= 308 ;
				WHEN  143  =>
					 sin_pos <= 311 ;
				WHEN  144  =>
					 sin_pos <= 314 ;
				WHEN  145  =>
					 sin_pos <= 317 ;
				WHEN  146  =>
					 sin_pos <= 320 ;
				WHEN  147  =>
					 sin_pos <= 323 ;
				WHEN  148  =>
					 sin_pos <= 326 ;
				WHEN  149  =>
					 sin_pos <= 328 ;
				WHEN  150  =>
					 sin_pos <= 331 ;
				WHEN  151  =>
					 sin_pos <= 334 ;
				WHEN  152  =>
					 sin_pos <= 337 ;
				WHEN  153  =>
					 sin_pos <= 340 ;
				WHEN  154  =>
					 sin_pos <= 343 ;
				WHEN  155  =>
					 sin_pos <= 346 ;
				WHEN  156  =>
					 sin_pos <= 348 ;
				WHEN  157  =>
					 sin_pos <= 351 ;
				WHEN  158  =>
					 sin_pos <= 354 ;
				WHEN  159  =>
					 sin_pos <= 357 ;
				WHEN  160  =>
					 sin_pos <= 359 ;
				WHEN  161  =>
					 sin_pos <= 362 ;
				WHEN  162  =>
					 sin_pos <= 365 ;
				WHEN  163  =>
					 sin_pos <= 368 ;
				WHEN  164  =>
					 sin_pos <= 370 ;
				WHEN  165  =>
					 sin_pos <= 373 ;
				WHEN  166  =>
					 sin_pos <= 375 ;
				WHEN  167  =>
					 sin_pos <= 378 ;
				WHEN  168  =>
					 sin_pos <= 381 ;
				WHEN  169  =>
					 sin_pos <= 383 ;
				WHEN  170  =>
					 sin_pos <= 386 ;
				WHEN  171  =>
					 sin_pos <= 388 ;
				WHEN  172  =>
					 sin_pos <= 391 ;
				WHEN  173  =>
					 sin_pos <= 393 ;
				WHEN  174  =>
					 sin_pos <= 395 ;
				WHEN  175  =>
					 sin_pos <= 398 ;
				WHEN  176  =>
					 sin_pos <= 400 ;
				WHEN  177  =>
					 sin_pos <= 402 ;
				WHEN  178  =>
					 sin_pos <= 405 ;
				WHEN  179  =>
					 sin_pos <= 407 ;
				WHEN  180  =>
					 sin_pos <= 409 ;
				WHEN  181  =>
					 sin_pos <= 411 ;
				WHEN  182  =>
					 sin_pos <= 414 ;
				WHEN  183  =>
					 sin_pos <= 416 ;
				WHEN  184  =>
					 sin_pos <= 418 ;
				WHEN  185  =>
					 sin_pos <= 420 ;
				WHEN  186  =>
					 sin_pos <= 422 ;
				WHEN  187  =>
					 sin_pos <= 424 ;
				WHEN  188  =>
					 sin_pos <= 426 ;
				WHEN  189  =>
					 sin_pos <= 428 ;
				WHEN  190  =>
					 sin_pos <= 430 ;
				WHEN  191  =>
					 sin_pos <= 432 ;
				WHEN  192  =>
					 sin_pos <= 434 ;
				WHEN  193  =>
					 sin_pos <= 435 ;
				WHEN  194  =>
					 sin_pos <= 437 ;
				WHEN  195  =>
					 sin_pos <= 439 ;
				WHEN  196  =>
					 sin_pos <= 441 ;
				WHEN  197  =>
					 sin_pos <= 442 ;
				WHEN  198  =>
					 sin_pos <= 444 ;
				WHEN  199  =>
					 sin_pos <= 446 ;
				WHEN  200  =>
					 sin_pos <= 447 ;
				WHEN  201  =>
					 sin_pos <= 449 ;
				WHEN  202  =>
					 sin_pos <= 450 ;
				WHEN  203  =>
					 sin_pos <= 452 ;
				WHEN  204  =>
					 sin_pos <= 453 ;
				WHEN  205  =>
					 sin_pos <= 455 ;
				WHEN  206  =>
					 sin_pos <= 456 ;
				WHEN  207  =>
					 sin_pos <= 457 ;
				WHEN  208  =>
					 sin_pos <= 459 ;
				WHEN  209  =>
					 sin_pos <= 460 ;
				WHEN  210  =>
					 sin_pos <= 461 ;
				WHEN  211  =>
					 sin_pos <= 462 ;
				WHEN  212  =>
					 sin_pos <= 464 ;
				WHEN  213  =>
					 sin_pos <= 465 ;
				WHEN  214  =>
					 sin_pos <= 466 ;
				WHEN  215  =>
					 sin_pos <= 467 ;
				WHEN  216  =>
					 sin_pos <= 468 ;
				WHEN  217  =>
					 sin_pos <= 469 ;
				WHEN  218  =>
					 sin_pos <= 470 ;
				WHEN  219  =>
					 sin_pos <= 470 ;
				WHEN  220  =>
					 sin_pos <= 471 ;
				WHEN  221  =>
					 sin_pos <= 472 ;
				WHEN  222  =>
					 sin_pos <= 473 ;
				WHEN  223  =>
					 sin_pos <= 474 ;
				WHEN  224  =>
					 sin_pos <= 474 ;
				WHEN  225  =>
					 sin_pos <= 475 ;
				WHEN  226  =>
					 sin_pos <= 475 ;
				WHEN  227  =>
					 sin_pos <= 476 ;
				WHEN  228  =>
					 sin_pos <= 477 ;
				WHEN  229  =>
					 sin_pos <= 477 ;
				WHEN  230  =>
					 sin_pos <= 477 ;
				WHEN  231  =>
					 sin_pos <= 478 ;
				WHEN  232  =>
					 sin_pos <= 478 ;
				WHEN  233  =>
					 sin_pos <= 478 ;
				WHEN  234  =>
					 sin_pos <= 479 ;
				WHEN  235  =>
					 sin_pos <= 479 ;
				WHEN  236  =>
					 sin_pos <= 479 ;
				WHEN  237  =>
					 sin_pos <= 479 ;
				WHEN  238  =>
					 sin_pos <= 479 ;
				WHEN  239  =>
					 sin_pos <= 479 ;
				WHEN  240  =>
					 sin_pos <= 479 ;
				WHEN  241  =>
					 sin_pos <= 479 ;
				WHEN  242  =>
					 sin_pos <= 479 ;
				WHEN  243  =>
					 sin_pos <= 479 ;
				WHEN  244  =>
					 sin_pos <= 479 ;
				WHEN  245  =>
					 sin_pos <= 479 ;
				WHEN  246  =>
					 sin_pos <= 479 ;
				WHEN  247  =>
					 sin_pos <= 478 ;
				WHEN  248  =>
					 sin_pos <= 478 ;
				WHEN  249  =>
					 sin_pos <= 478 ;
				WHEN  250  =>
					 sin_pos <= 477 ;
				WHEN  251  =>
					 sin_pos <= 477 ;
				WHEN  252  =>
					 sin_pos <= 477 ;
				WHEN  253  =>
					 sin_pos <= 476 ;
				WHEN  254  =>
					 sin_pos <= 475 ;
				WHEN  255  =>
					 sin_pos <= 475 ;
				WHEN  256  =>
					 sin_pos <= 474 ;
				WHEN  257  =>
					 sin_pos <= 474 ;
				WHEN  258  =>
					 sin_pos <= 473 ;
				WHEN  259  =>
					 sin_pos <= 472 ;
				WHEN  260  =>
					 sin_pos <= 471 ;
				WHEN  261  =>
					 sin_pos <= 470 ;
				WHEN  262  =>
					 sin_pos <= 470 ;
				WHEN  263  =>
					 sin_pos <= 469 ;
				WHEN  264  =>
					 sin_pos <= 468 ;
				WHEN  265  =>
					 sin_pos <= 467 ;
				WHEN  266  =>
					 sin_pos <= 466 ;
				WHEN  267  =>
					 sin_pos <= 465 ;
				WHEN  268  =>
					 sin_pos <= 464 ;
				WHEN  269  =>
					 sin_pos <= 462 ;
				WHEN  270  =>
					 sin_pos <= 461 ;
				WHEN  271  =>
					 sin_pos <= 460 ;
				WHEN  272  =>
					 sin_pos <= 459 ;
				WHEN  273  =>
					 sin_pos <= 457 ;
				WHEN  274  =>
					 sin_pos <= 456 ;
				WHEN  275  =>
					 sin_pos <= 455 ;
				WHEN  276  =>
					 sin_pos <= 453 ;
				WHEN  277  =>
					 sin_pos <= 452 ;
				WHEN  278  =>
					 sin_pos <= 450 ;
				WHEN  279  =>
					 sin_pos <= 449 ;
				WHEN  280  =>
					 sin_pos <= 447 ;
				WHEN  281  =>
					 sin_pos <= 446 ;
				WHEN  282  =>
					 sin_pos <= 444 ;
				WHEN  283  =>
					 sin_pos <= 442 ;
				WHEN  284  =>
					 sin_pos <= 441 ;
				WHEN  285  =>
					 sin_pos <= 439 ;
				WHEN  286  =>
					 sin_pos <= 437 ;
				WHEN  287  =>
					 sin_pos <= 435 ;
				WHEN  288  =>
					 sin_pos <= 434 ;
				WHEN  289  =>
					 sin_pos <= 432 ;
				WHEN  290  =>
					 sin_pos <= 430 ;
				WHEN  291  =>
					 sin_pos <= 428 ;
				WHEN  292  =>
					 sin_pos <= 426 ;
				WHEN  293  =>
					 sin_pos <= 424 ;
				WHEN  294  =>
					 sin_pos <= 422 ;
				WHEN  295  =>
					 sin_pos <= 420 ;
				WHEN  296  =>
					 sin_pos <= 418 ;
				WHEN  297  =>
					 sin_pos <= 416 ;
				WHEN  298  =>
					 sin_pos <= 414 ;
				WHEN  299  =>
					 sin_pos <= 411 ;
				WHEN  300  =>
					 sin_pos <= 409 ;
				WHEN  301  =>
					 sin_pos <= 407 ;
				WHEN  302  =>
					 sin_pos <= 405 ;
				WHEN  303  =>
					 sin_pos <= 402 ;
				WHEN  304  =>
					 sin_pos <= 400 ;
				WHEN  305  =>
					 sin_pos <= 398 ;
				WHEN  306  =>
					 sin_pos <= 395 ;
				WHEN  307  =>
					 sin_pos <= 393 ;
				WHEN  308  =>
					 sin_pos <= 391 ;
				WHEN  309  =>
					 sin_pos <= 388 ;
				WHEN  310  =>
					 sin_pos <= 386 ;
				WHEN  311  =>
					 sin_pos <= 383 ;
				WHEN  312  =>
					 sin_pos <= 381 ;
				WHEN  313  =>
					 sin_pos <= 378 ;
				WHEN  314  =>
					 sin_pos <= 375 ;
				WHEN  315  =>
					 sin_pos <= 373 ;
				WHEN  316  =>
					 sin_pos <= 370 ;
				WHEN  317  =>
					 sin_pos <= 368 ;
				WHEN  318  =>
					 sin_pos <= 365 ;
				WHEN  319  =>
					 sin_pos <= 362 ;
				WHEN  320  =>
					 sin_pos <= 360 ;
				WHEN  321  =>
					 sin_pos <= 357 ;
				WHEN  322  =>
					 sin_pos <= 354 ;
				WHEN  323  =>
					 sin_pos <= 351 ;
				WHEN  324  =>
					 sin_pos <= 348 ;
				WHEN  325  =>
					 sin_pos <= 346 ;
				WHEN  326  =>
					 sin_pos <= 343 ;
				WHEN  327  =>
					 sin_pos <= 340 ;
				WHEN  328  =>
					 sin_pos <= 337 ;
				WHEN  329  =>
					 sin_pos <= 334 ;
				WHEN  330  =>
					 sin_pos <= 331 ;
				WHEN  331  =>
					 sin_pos <= 328 ;
				WHEN  332  =>
					 sin_pos <= 326 ;
				WHEN  333  =>
					 sin_pos <= 323 ;
				WHEN  334  =>
					 sin_pos <= 320 ;
				WHEN  335  =>
					 sin_pos <= 317 ;
				WHEN  336  =>
					 sin_pos <= 314 ;
				WHEN  337  =>
					 sin_pos <= 311 ;
				WHEN  338  =>
					 sin_pos <= 308 ;
				WHEN  339  =>
					 sin_pos <= 305 ;
				WHEN  340  =>
					 sin_pos <= 302 ;
				WHEN  341  =>
					 sin_pos <= 299 ;
				WHEN  342  =>
					 sin_pos <= 296 ;
				WHEN  343  =>
					 sin_pos <= 292 ;
				WHEN  344  =>
					 sin_pos <= 289 ;
				WHEN  345  =>
					 sin_pos <= 286 ;
				WHEN  346  =>
					 sin_pos <= 283 ;
				WHEN  347  =>
					 sin_pos <= 280 ;
				WHEN  348  =>
					 sin_pos <= 277 ;
				WHEN  349  =>
					 sin_pos <= 274 ;
				WHEN  350  =>
					 sin_pos <= 271 ;
				WHEN  351  =>
					 sin_pos <= 268 ;
				WHEN  352  =>
					 sin_pos <= 265 ;
				WHEN  353  =>
					 sin_pos <= 261 ;
				WHEN  354  =>
					 sin_pos <= 258 ;
				WHEN  355  =>
					 sin_pos <= 255 ;
				WHEN  356  =>
					 sin_pos <= 252 ;
				WHEN  357  =>
					 sin_pos <= 249 ;
				WHEN  358  =>
					 sin_pos <= 246 ;
				WHEN  359  =>
					 sin_pos <= 243 ;
				WHEN  360  =>
					 sin_pos <= 240 ;
				WHEN  361  =>
					 sin_pos <= 236 ;
				WHEN  362  =>
					 sin_pos <= 233 ;
				WHEN  363  =>
					 sin_pos <= 230 ;
				WHEN  364  =>
					 sin_pos <= 227 ;
				WHEN  365  =>
					 sin_pos <= 224 ;
				WHEN  366  =>
					 sin_pos <= 221 ;
				WHEN  367  =>
					 sin_pos <= 218 ;
				WHEN  368  =>
					 sin_pos <= 214 ;
				WHEN  369  =>
					 sin_pos <= 211 ;
				WHEN  370  =>
					 sin_pos <= 208 ;
				WHEN  371  =>
					 sin_pos <= 205 ;
				WHEN  372  =>
					 sin_pos <= 202 ;
				WHEN  373  =>
					 sin_pos <= 199 ;
				WHEN  374  =>
					 sin_pos <= 196 ;
				WHEN  375  =>
					 sin_pos <= 193 ;
				WHEN  376  =>
					 sin_pos <= 190 ;
				WHEN  377  =>
					 sin_pos <= 187 ;
				WHEN  378  =>
					 sin_pos <= 183 ;
				WHEN  379  =>
					 sin_pos <= 180 ;
				WHEN  380  =>
					 sin_pos <= 177 ;
				WHEN  381  =>
					 sin_pos <= 174 ;
				WHEN  382  =>
					 sin_pos <= 171 ;
				WHEN  383  =>
					 sin_pos <= 168 ;
				WHEN  384  =>
					 sin_pos <= 165 ;
				WHEN  385  =>
					 sin_pos <= 162 ;
				WHEN  386  =>
					 sin_pos <= 159 ;
				WHEN  387  =>
					 sin_pos <= 156 ;
				WHEN  388  =>
					 sin_pos <= 153 ;
				WHEN  389  =>
					 sin_pos <= 151 ;
				WHEN  390  =>
					 sin_pos <= 148 ;
				WHEN  391  =>
					 sin_pos <= 145 ;
				WHEN  392  =>
					 sin_pos <= 142 ;
				WHEN  393  =>
					 sin_pos <= 139 ;
				WHEN  394  =>
					 sin_pos <= 136 ;
				WHEN  395  =>
					 sin_pos <= 133 ;
				WHEN  396  =>
					 sin_pos <= 131 ;
				WHEN  397  =>
					 sin_pos <= 128 ;
				WHEN  398  =>
					 sin_pos <= 125 ;
				WHEN  399  =>
					 sin_pos <= 122 ;
				WHEN  400  =>
					 sin_pos <= 119 ;
				WHEN  401  =>
					 sin_pos <= 117 ;
				WHEN  402  =>
					 sin_pos <= 114 ;
				WHEN  403  =>
					 sin_pos <= 111 ;
				WHEN  404  =>
					 sin_pos <= 109 ;
				WHEN  405  =>
					 sin_pos <= 106 ;
				WHEN  406  =>
					 sin_pos <= 104 ;
				WHEN  407  =>
					 sin_pos <= 101 ;
				WHEN  408  =>
					 sin_pos <= 98 ;
				WHEN  409  =>
					 sin_pos <= 96 ;
				WHEN  410  =>
					 sin_pos <= 93 ;
				WHEN  411  =>
					 sin_pos <= 91 ;
				WHEN  412  =>
					 sin_pos <= 88 ;
				WHEN  413  =>
					 sin_pos <= 86 ;
				WHEN  414  =>
					 sin_pos <= 84 ;
				WHEN  415  =>
					 sin_pos <= 81 ;
				WHEN  416  =>
					 sin_pos <= 79 ;
				WHEN  417  =>
					 sin_pos <= 77 ;
				WHEN  418  =>
					 sin_pos <= 74 ;
				WHEN  419  =>
					 sin_pos <= 72 ;
				WHEN  420  =>
					 sin_pos <= 70 ;
				WHEN  421  =>
					 sin_pos <= 68 ;
				WHEN  422  =>
					 sin_pos <= 65 ;
				WHEN  423  =>
					 sin_pos <= 63 ;
				WHEN  424  =>
					 sin_pos <= 61 ;
				WHEN  425  =>
					 sin_pos <= 59 ;
				WHEN  426  =>
					 sin_pos <= 57 ;
				WHEN  427  =>
					 sin_pos <= 55 ;
				WHEN  428  =>
					 sin_pos <= 53 ;
				WHEN  429  =>
					 sin_pos <= 51 ;
				WHEN  430  =>
					 sin_pos <= 49 ;
				WHEN  431  =>
					 sin_pos <= 47 ;
				WHEN  432  =>
					 sin_pos <= 45 ;
				WHEN  433  =>
					 sin_pos <= 44 ;
				WHEN  434  =>
					 sin_pos <= 42 ;
				WHEN  435  =>
					 sin_pos <= 40 ;
				WHEN  436  =>
					 sin_pos <= 38 ;
				WHEN  437  =>
					 sin_pos <= 37 ;
				WHEN  438  =>
					 sin_pos <= 35 ;
				WHEN  439  =>
					 sin_pos <= 33 ;
				WHEN  440  =>
					 sin_pos <= 32 ;
				WHEN  441  =>
					 sin_pos <= 30 ;
				WHEN  442  =>
					 sin_pos <= 29 ;
				WHEN  443  =>
					 sin_pos <= 27 ;
				WHEN  444  =>
					 sin_pos <= 26 ;
				WHEN  445  =>
					 sin_pos <= 24 ;
				WHEN  446  =>
					 sin_pos <= 23 ;
				WHEN  447  =>
					 sin_pos <= 22 ;
				WHEN  448  =>
					 sin_pos <= 20 ;
				WHEN  449  =>
					 sin_pos <= 19 ;
				WHEN  450  =>
					 sin_pos <= 18 ;
				WHEN  451  =>
					 sin_pos <= 17 ;
				WHEN  452  =>
					 sin_pos <= 15 ;
				WHEN  453  =>
					 sin_pos <= 14 ;
				WHEN  454  =>
					 sin_pos <= 13 ;
				WHEN  455  =>
					 sin_pos <= 12 ;
				WHEN  456  =>
					 sin_pos <= 11 ;
				WHEN  457  =>
					 sin_pos <= 10 ;
				WHEN  458  =>
					 sin_pos <= 9 ;
				WHEN  459  =>
					 sin_pos <= 9 ;
				WHEN  460  =>
					 sin_pos <= 8 ;
				WHEN  461  =>
					 sin_pos <= 7 ;
				WHEN  462  =>
					 sin_pos <= 6 ;
				WHEN  463  =>
					 sin_pos <= 5 ;
				WHEN  464  =>
					 sin_pos <= 5 ;
				WHEN  465  =>
					 sin_pos <= 4 ;
				WHEN  466  =>
					 sin_pos <= 4 ;
				WHEN  467  =>
					 sin_pos <= 3 ;
				WHEN  468  =>
					 sin_pos <= 2 ;
				WHEN  469  =>
					 sin_pos <= 2 ;
				WHEN  470  =>
					 sin_pos <= 2 ;
				WHEN  471  =>
					 sin_pos <= 1 ;
				WHEN  472  =>
					 sin_pos <= 1 ;
				WHEN  473  =>
					 sin_pos <= 1 ;
				WHEN  474  =>
					 sin_pos <= 0 ;
				WHEN  475  =>
					 sin_pos <= 0 ;
				WHEN  476  =>
					 sin_pos <= 0 ;
				WHEN  477  =>
					 sin_pos <= 0 ;
				WHEN  478  =>
					 sin_pos <= 0 ;
				WHEN  479  =>
					 sin_pos <= 0 ;
				WHEN OTHERS =>	 
					sin_pos <= 0;
			END CASE;
			
			Delay_reg(0) <= In1_signed;
			Delay_reg(1 TO 479) <= Delay_reg(0 TO 478);
      END IF;
    END IF;
  END PROCESS Delay_process;

  Delay_out1 <= Delay_reg(sin_pos);

  attenuation_cast <= resize(Delay_out1 & '0' & '0' & '0' & '0' & '0' & '0', 16);
  attenuation_out1 <= attenuation_cast(14 DOWNTO 7) + ('0' & (attenuation_cast(6) AND (( NOT attenuation_cast(15)) OR (attenuation_cast(5) OR attenuation_cast(4) OR attenuation_cast(3) OR attenuation_cast(2) OR attenuation_cast(1) OR attenuation_cast(0)))));
  attenuation_cast2 <= resize(In1_signed & '0' & '0' & '0' & '0' & '0' & '0', 16);
  attenuation_out2 <= attenuation_cast2(14 DOWNTO 7) + ('0' & (attenuation_cast2(6) AND (( NOT attenuation_cast2(15)) OR (attenuation_cast2(5) OR attenuation_cast2(4) OR attenuation_cast2(3) OR attenuation_cast2(2) OR attenuation_cast2(1) OR attenuation_cast2(0)))));
  Sum_out1 <= attenuation_out2 + attenuation_out1;

  Out1 <= std_logic_vector(Sum_out1);

  ce_out <= clk_enable;

END rtl;
